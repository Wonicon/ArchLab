module misp_cpu_top (
    input clk
);

reg [31:0] PC;


endmodule
